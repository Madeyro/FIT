-- fsm.vhd: Finite State Machine
-- Author(s): Maros Kopec, xkopec44
-- kod1 = 1245164665     kod2 = 12451675984

library ieee;
use ieee.std_logic_1164.all;
-- ----------------------------------------------------------------------------
--                        Entity declaration
-- ----------------------------------------------------------------------------
entity fsm is
port(
   CLK         : in  std_logic;
   RESET       : in  std_logic;

   -- Input signals
   KEY         : in  std_logic_vector(15 downto 0);
   CNT_OF      : in  std_logic;

   -- Output signals
   FSM_CNT_CE  : out std_logic;
   FSM_MX_MEM  : out std_logic;
   FSM_MX_LCD  : out std_logic;
   FSM_LCD_WR  : out std_logic;
   FSM_LCD_CLR : out std_logic
);
end entity fsm;

-- ----------------------------------------------------------------------------
--                      Architecture declaration
-- ----------------------------------------------------------------------------
architecture behavioral of fsm is
   type t_state is (FAIL, TEST_NO1, TEST_NO2, TEST_NO3, TEST_NO4, TEST_NO5,
                     TEST_NO6, TEST_NO7, TEST_NO8A, TEST_NO8B, TEST_NO9A, TEST_NO9B,
                     TEST_NO10A, TEST_NO10B, TEST_NO11, TEST_CNF,
                     PRINT_FAILED, PRINT_SUCCESSFUL, FINISH);
   signal present_state, next_state : t_state;

begin
-- -------------------------------------------------------
sync_logic : process(RESET, CLK)
begin
   if (RESET = '1') then
      present_state <= TEST_NO1;
   elsif (CLK'event AND CLK = '1') then
      present_state <= next_state;
   end if;
end process sync_logic;

-- -------------------------------------------------------
next_state_logic : process(present_state, KEY, CNT_OF)
begin
   case (present_state) is
   -- --------------------------------------------
   when FAIL =>
      next_state <= FAIL;
      if (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO1 =>
      next_state <= TEST_NO1;
      if (KEY(1) = '1') then
         next_state <= TEST_NO2; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO2 =>
      next_state <= TEST_NO2;
      if (KEY(2) = '1') then
         next_state <= TEST_NO3; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO3 =>
      next_state <= TEST_NO3;
      if (KEY(4) = '1') then
         next_state <= TEST_NO4; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO4 =>
      next_state <= TEST_NO4;
      if (KEY(5) = '1') then
         next_state <= TEST_NO5; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO5 =>
      next_state <= TEST_NO5;
      if (KEY(1) = '1') then
         next_state <= TEST_NO6; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO6 =>
      next_state <= TEST_NO6;
      if (KEY(6) = '1') then
         next_state <= TEST_NO7; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO7 =>
      next_state <= TEST_NO7;
      if (KEY(4) = '1') then
         next_state <= TEST_NO8A;
      elsif (KEY(7) = '1') then
         next_state <= TEST_NO8B;
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO8A =>
      next_state <= TEST_NO8A;
      if (KEY(6) = '1') then
         next_state <= TEST_NO9A; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO8B =>
      next_state <= TEST_NO8B;
      if (KEY(5) = '1') then
         next_state <= TEST_NO9B; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO9A =>
      next_state <= TEST_NO9A;
      if (KEY(6) = '1') then
         next_state <= TEST_NO10A; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO9B =>
      next_state <= TEST_NO9B;
      if (KEY(9) = '1') then
         next_state <= TEST_NO10B; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO10A =>
      next_state <= TEST_NO10A;
      if (KEY(5) = '1') then
         next_state <= TEST_CNF; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO10B =>
      next_state <= TEST_NO10B;
      if (KEY(8) = '1') then
         next_state <= TEST_NO11; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_NO11 =>
      next_state <= TEST_NO11;
      if (KEY(4) = '1') then
         next_state <= TEST_CNF; 
      elsif (KEY(15) = '1') then
         next_state <= PRINT_FAILED;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
      -- - - - - - - - - - - - - - - - - - - - - - -
   when TEST_CNF =>
      next_state <= TEST_CNF;
      if (KEY(15) = '1') then
         next_state <= PRINT_SUCCESSFUL;
      elsif (KEY(15 downto 0) /= "0000000000000000") then
         next_state <= FAIL;
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when PRINT_SUCCESSFUL => 
      next_state <= PRINT_SUCCESSFUL;
      if (CNT_OF = '1') then
         next_state <= FINISH;
      end if;
      -- --------------------------------------------
   when PRINT_FAILED =>
      next_state <= PRINT_FAILED;
      if (CNT_OF = '1') then
         next_state <= FINISH;
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when FINISH =>
      next_state <= FINISH;
      if (KEY(15) = '1') then
         next_state <= TEST_NO1; 
      end if;
   -- - - - - - - - - - - - - - - - - - - - - - -
   when others =>
      next_state <= TEST_NO1;
   end case;
end process next_state_logic;

-- -------------------------------------------------------
output_logic : process(present_state, KEY)
begin
   FSM_CNT_CE     <= '0';
   FSM_MX_MEM     <= '0';
   FSM_MX_LCD     <= '0';
   FSM_LCD_WR     <= '0';
   FSM_LCD_CLR    <= '0';

   case (present_state) is
   -- - - - - - - - - - - - - - - - - - - - - - -
   when PRINT_FAILED =>
      FSM_CNT_CE     <= '1';
      FSM_MX_LCD     <= '1';
      FSM_MX_MEM     <= '0';
      FSM_LCD_WR     <= '1';
 
   -- - - - - - - - - - - - - - - - - - - - - - -
   when PRINT_SUCCESSFUL =>
      FSM_CNT_CE     <= '1';
      FSM_MX_LCD     <= '1';
      FSM_MX_MEM     <= '1';
      FSM_LCD_WR     <= '1';
 
   -- - - - - - - - - - - - - - - - - - - - - - -
   when FINISH =>
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
 
   -- - - - - - - - - - - - - - - - - - - - - - -
   when others =>
   if (KEY(14 downto 0) /= "000000000000000") then
         FSM_LCD_WR     <= '1';
      end if;
      if (KEY(15) = '1') then
         FSM_LCD_CLR    <= '1';
      end if;
   end case;
end process output_logic;
 
end architecture behavioral;